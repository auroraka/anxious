// anxious_qsys_tb.v

// Generated using ACDS version 15.0 145

`timescale 1 ns / 1 ns
module anxious_qsys_tb (
	);

	wire         anxious_qsys_inst_clk_bfm_clk_clk;                            // anxious_qsys_inst_clk_bfm:clk -> [anxious_qsys_inst:clk_clk, anxious_qsys_inst_reset_bfm:clk]
	wire         sdram_controller_0_my_partner_clk_bfm_clk_clk;                // sdram_controller_0_my_partner_clk_bfm:clk -> sdram_controller_0_my_partner:clk
	wire   [0:0] anxious_qsys_inst_camera_mm_0_conduit_bfm_conduit_cam_vsync;  // anxious_qsys_inst_camera_mm_0_conduit_bfm:sig_cam_vsync -> anxious_qsys_inst:camera_mm_0_conduit_cam_vsync
	wire         anxious_qsys_inst_camera_mm_0_conduit_cam_pwdn;               // anxious_qsys_inst:camera_mm_0_conduit_cam_pwdn -> anxious_qsys_inst_camera_mm_0_conduit_bfm:sig_cam_pwdn
	wire   [7:0] anxious_qsys_inst_camera_mm_0_conduit_bfm_conduit_cam_din;    // anxious_qsys_inst_camera_mm_0_conduit_bfm:sig_cam_din -> anxious_qsys_inst:camera_mm_0_conduit_cam_din
	wire   [0:0] anxious_qsys_inst_camera_mm_0_conduit_bfm_conduit_cam_pclk;   // anxious_qsys_inst_camera_mm_0_conduit_bfm:sig_cam_pclk -> anxious_qsys_inst:camera_mm_0_conduit_cam_pclk
	wire   [0:0] anxious_qsys_inst_camera_mm_0_conduit_bfm_conduit_enable_n;   // anxious_qsys_inst_camera_mm_0_conduit_bfm:sig_enable_n -> anxious_qsys_inst:camera_mm_0_conduit_enable_n
	wire   [0:0] anxious_qsys_inst_camera_mm_0_conduit_bfm_conduit_cam_href;   // anxious_qsys_inst_camera_mm_0_conduit_bfm:sig_cam_href -> anxious_qsys_inst:camera_mm_0_conduit_cam_href
	wire         anxious_qsys_inst_camera_mm_0_conduit_cam_xclk;               // anxious_qsys_inst:camera_mm_0_conduit_cam_xclk -> anxious_qsys_inst_camera_mm_0_conduit_bfm:sig_cam_xclk
	wire         anxious_qsys_inst_camera_mm_0_conduit_cam_reset;              // anxious_qsys_inst:camera_mm_0_conduit_cam_reset -> anxious_qsys_inst_camera_mm_0_conduit_bfm:sig_cam_reset
	wire   [0:0] anxious_qsys_inst_camera_mm_0_conduit_bfm_conduit_clk_camera; // anxious_qsys_inst_camera_mm_0_conduit_bfm:sig_clk_camera -> anxious_qsys_inst:camera_mm_0_conduit_clk_camera
	wire   [7:0] anxious_qsys_inst_led_export;                                 // anxious_qsys_inst:led_export -> anxious_qsys_inst_led_bfm:sig_export
	wire         anxious_qsys_inst_new_sdram_controller_0_wire_cs_n;           // anxious_qsys_inst:new_sdram_controller_0_wire_cs_n -> sdram_controller_0_my_partner:zs_cs_n
	wire   [3:0] anxious_qsys_inst_new_sdram_controller_0_wire_dqm;            // anxious_qsys_inst:new_sdram_controller_0_wire_dqm -> sdram_controller_0_my_partner:zs_dqm
	wire         anxious_qsys_inst_new_sdram_controller_0_wire_cas_n;          // anxious_qsys_inst:new_sdram_controller_0_wire_cas_n -> sdram_controller_0_my_partner:zs_cas_n
	wire         anxious_qsys_inst_new_sdram_controller_0_wire_ras_n;          // anxious_qsys_inst:new_sdram_controller_0_wire_ras_n -> sdram_controller_0_my_partner:zs_ras_n
	wire         anxious_qsys_inst_new_sdram_controller_0_wire_we_n;           // anxious_qsys_inst:new_sdram_controller_0_wire_we_n -> sdram_controller_0_my_partner:zs_we_n
	wire  [12:0] anxious_qsys_inst_new_sdram_controller_0_wire_addr;           // anxious_qsys_inst:new_sdram_controller_0_wire_addr -> sdram_controller_0_my_partner:zs_addr
	wire         anxious_qsys_inst_new_sdram_controller_0_wire_cke;            // anxious_qsys_inst:new_sdram_controller_0_wire_cke -> sdram_controller_0_my_partner:zs_cke
	wire  [31:0] anxious_qsys_inst_new_sdram_controller_0_wire_dq;             // [] -> [anxious_qsys_inst:new_sdram_controller_0_wire_dq, sdram_controller_0_my_partner:zs_dq]
	wire   [1:0] anxious_qsys_inst_new_sdram_controller_0_wire_ba;             // anxious_qsys_inst:new_sdram_controller_0_wire_ba -> sdram_controller_0_my_partner:zs_ba
	wire         anxious_qsys_inst_vga_mm_0_conduit_vga_clk;                   // anxious_qsys_inst:vga_mm_0_conduit_vga_clk -> anxious_qsys_inst_vga_mm_0_conduit_bfm:sig_vga_clk
	wire   [0:0] anxious_qsys_inst_vga_mm_0_conduit_bfm_conduit_clk_vga;       // anxious_qsys_inst_vga_mm_0_conduit_bfm:sig_clk_vga -> anxious_qsys_inst:vga_mm_0_conduit_clk_vga
	wire   [7:0] anxious_qsys_inst_vga_mm_0_conduit_vga_g;                     // anxious_qsys_inst:vga_mm_0_conduit_vga_g -> anxious_qsys_inst_vga_mm_0_conduit_bfm:sig_vga_g
	wire         anxious_qsys_inst_vga_mm_0_conduit_vga_sync_n;                // anxious_qsys_inst:vga_mm_0_conduit_vga_sync_n -> anxious_qsys_inst_vga_mm_0_conduit_bfm:sig_vga_sync_n
	wire         anxious_qsys_inst_vga_mm_0_conduit_vga_vs;                    // anxious_qsys_inst:vga_mm_0_conduit_vga_vs -> anxious_qsys_inst_vga_mm_0_conduit_bfm:sig_vga_vs
	wire         anxious_qsys_inst_vga_mm_0_conduit_vga_blank_n;               // anxious_qsys_inst:vga_mm_0_conduit_vga_blank_n -> anxious_qsys_inst_vga_mm_0_conduit_bfm:sig_vga_blank_n
	wire   [7:0] anxious_qsys_inst_vga_mm_0_conduit_vga_b;                     // anxious_qsys_inst:vga_mm_0_conduit_vga_b -> anxious_qsys_inst_vga_mm_0_conduit_bfm:sig_vga_b
	wire   [7:0] anxious_qsys_inst_vga_mm_0_conduit_vga_r;                     // anxious_qsys_inst:vga_mm_0_conduit_vga_r -> anxious_qsys_inst_vga_mm_0_conduit_bfm:sig_vga_r
	wire         anxious_qsys_inst_vga_mm_0_conduit_vga_hs;                    // anxious_qsys_inst:vga_mm_0_conduit_vga_hs -> anxious_qsys_inst_vga_mm_0_conduit_bfm:sig_vga_hs
	wire         anxious_qsys_inst_reset_bfm_reset_reset;                      // anxious_qsys_inst_reset_bfm:reset -> anxious_qsys_inst:reset_reset_n

	anxious_qsys anxious_qsys_inst (
		.camera_mm_0_conduit_clk_camera    (anxious_qsys_inst_camera_mm_0_conduit_bfm_conduit_clk_camera), //         camera_mm_0_conduit.clk_camera
		.camera_mm_0_conduit_enable_n      (anxious_qsys_inst_camera_mm_0_conduit_bfm_conduit_enable_n),   //                            .enable_n
		.camera_mm_0_conduit_cam_din       (anxious_qsys_inst_camera_mm_0_conduit_bfm_conduit_cam_din),    //                            .cam_din
		.camera_mm_0_conduit_cam_href      (anxious_qsys_inst_camera_mm_0_conduit_bfm_conduit_cam_href),   //                            .cam_href
		.camera_mm_0_conduit_cam_pclk      (anxious_qsys_inst_camera_mm_0_conduit_bfm_conduit_cam_pclk),   //                            .cam_pclk
		.camera_mm_0_conduit_cam_pwdn      (anxious_qsys_inst_camera_mm_0_conduit_cam_pwdn),               //                            .cam_pwdn
		.camera_mm_0_conduit_cam_reset     (anxious_qsys_inst_camera_mm_0_conduit_cam_reset),              //                            .cam_reset
		.camera_mm_0_conduit_cam_vsync     (anxious_qsys_inst_camera_mm_0_conduit_bfm_conduit_cam_vsync),  //                            .cam_vsync
		.camera_mm_0_conduit_cam_xclk      (anxious_qsys_inst_camera_mm_0_conduit_cam_xclk),               //                            .cam_xclk
		.clk_clk                           (anxious_qsys_inst_clk_bfm_clk_clk),                            //                         clk.clk
		.led_export                        (anxious_qsys_inst_led_export),                                 //                         led.export
		.new_sdram_controller_0_wire_addr  (anxious_qsys_inst_new_sdram_controller_0_wire_addr),           // new_sdram_controller_0_wire.addr
		.new_sdram_controller_0_wire_ba    (anxious_qsys_inst_new_sdram_controller_0_wire_ba),             //                            .ba
		.new_sdram_controller_0_wire_cas_n (anxious_qsys_inst_new_sdram_controller_0_wire_cas_n),          //                            .cas_n
		.new_sdram_controller_0_wire_cke   (anxious_qsys_inst_new_sdram_controller_0_wire_cke),            //                            .cke
		.new_sdram_controller_0_wire_cs_n  (anxious_qsys_inst_new_sdram_controller_0_wire_cs_n),           //                            .cs_n
		.new_sdram_controller_0_wire_dq    (anxious_qsys_inst_new_sdram_controller_0_wire_dq),             //                            .dq
		.new_sdram_controller_0_wire_dqm   (anxious_qsys_inst_new_sdram_controller_0_wire_dqm),            //                            .dqm
		.new_sdram_controller_0_wire_ras_n (anxious_qsys_inst_new_sdram_controller_0_wire_ras_n),          //                            .ras_n
		.new_sdram_controller_0_wire_we_n  (anxious_qsys_inst_new_sdram_controller_0_wire_we_n),           //                            .we_n
		.reset_reset_n                     (anxious_qsys_inst_reset_bfm_reset_reset),                      //                       reset.reset_n
		.sys_sdram_pll_0_sdram_clk_clk     (),                                                             //   sys_sdram_pll_0_sdram_clk.clk
		.vga_mm_0_conduit_vga_b            (anxious_qsys_inst_vga_mm_0_conduit_vga_b),                     //            vga_mm_0_conduit.vga_b
		.vga_mm_0_conduit_vga_blank_n      (anxious_qsys_inst_vga_mm_0_conduit_vga_blank_n),               //                            .vga_blank_n
		.vga_mm_0_conduit_vga_clk          (anxious_qsys_inst_vga_mm_0_conduit_vga_clk),                   //                            .vga_clk
		.vga_mm_0_conduit_vga_g            (anxious_qsys_inst_vga_mm_0_conduit_vga_g),                     //                            .vga_g
		.vga_mm_0_conduit_vga_hs           (anxious_qsys_inst_vga_mm_0_conduit_vga_hs),                    //                            .vga_hs
		.vga_mm_0_conduit_vga_r            (anxious_qsys_inst_vga_mm_0_conduit_vga_r),                     //                            .vga_r
		.vga_mm_0_conduit_vga_sync_n       (anxious_qsys_inst_vga_mm_0_conduit_vga_sync_n),                //                            .vga_sync_n
		.vga_mm_0_conduit_vga_vs           (anxious_qsys_inst_vga_mm_0_conduit_vga_vs),                    //                            .vga_vs
		.vga_mm_0_conduit_clk_vga          (anxious_qsys_inst_vga_mm_0_conduit_bfm_conduit_clk_vga)        //                            .clk_vga
	);

	altera_conduit_bfm camera_bfm (
		.sig_clk_camera (anxious_qsys_inst_camera_mm_0_conduit_bfm_conduit_clk_camera), // conduit.clk_camera
		.sig_enable_n   (anxious_qsys_inst_camera_mm_0_conduit_bfm_conduit_enable_n),   //        .enable_n
		.sig_cam_din    (anxious_qsys_inst_camera_mm_0_conduit_bfm_conduit_cam_din),    //        .cam_din
		.sig_cam_href   (anxious_qsys_inst_camera_mm_0_conduit_bfm_conduit_cam_href),   //        .cam_href
		.sig_cam_pclk   (anxious_qsys_inst_camera_mm_0_conduit_bfm_conduit_cam_pclk),   //        .cam_pclk
		.sig_cam_pwdn   (anxious_qsys_inst_camera_mm_0_conduit_cam_pwdn),               //        .cam_pwdn
		.sig_cam_reset  (anxious_qsys_inst_camera_mm_0_conduit_cam_reset),              //        .cam_reset
		.sig_cam_vsync  (anxious_qsys_inst_camera_mm_0_conduit_bfm_conduit_cam_vsync),  //        .cam_vsync
		.sig_cam_xclk   (anxious_qsys_inst_camera_mm_0_conduit_cam_xclk)                //        .cam_xclk
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) anxious_qsys_inst_clk_bfm (
		.clk (anxious_qsys_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm_0002 anxious_qsys_inst_led_bfm (
		.sig_export (anxious_qsys_inst_led_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (6000)
	) anxious_qsys_inst_reset_bfm (
		.reset (anxious_qsys_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (anxious_qsys_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm_0003 anxious_qsys_inst_vga_mm_0_conduit_bfm (
		.sig_vga_b       (anxious_qsys_inst_vga_mm_0_conduit_vga_b),               // conduit.vga_b
		.sig_vga_blank_n (anxious_qsys_inst_vga_mm_0_conduit_vga_blank_n),         //        .vga_blank_n
		.sig_vga_clk     (anxious_qsys_inst_vga_mm_0_conduit_vga_clk),             //        .vga_clk
		.sig_vga_g       (anxious_qsys_inst_vga_mm_0_conduit_vga_g),               //        .vga_g
		.sig_vga_hs      (anxious_qsys_inst_vga_mm_0_conduit_vga_hs),              //        .vga_hs
		.sig_vga_r       (anxious_qsys_inst_vga_mm_0_conduit_vga_r),               //        .vga_r
		.sig_vga_sync_n  (anxious_qsys_inst_vga_mm_0_conduit_vga_sync_n),          //        .vga_sync_n
		.sig_vga_vs      (anxious_qsys_inst_vga_mm_0_conduit_vga_vs),              //        .vga_vs
		.sig_clk_vga     (anxious_qsys_inst_vga_mm_0_conduit_bfm_conduit_clk_vga)  //        .clk_vga
	);

	altera_sdram_partner_module sdram_controller_0_my_partner (
		.clk      (sdram_controller_0_my_partner_clk_bfm_clk_clk),       //     clk.clk
		.zs_dq    (anxious_qsys_inst_new_sdram_controller_0_wire_dq),    // conduit.dq
		.zs_addr  (anxious_qsys_inst_new_sdram_controller_0_wire_addr),  //        .addr
		.zs_ba    (anxious_qsys_inst_new_sdram_controller_0_wire_ba),    //        .ba
		.zs_cas_n (anxious_qsys_inst_new_sdram_controller_0_wire_cas_n), //        .cas_n
		.zs_cke   (anxious_qsys_inst_new_sdram_controller_0_wire_cke),   //        .cke
		.zs_cs_n  (anxious_qsys_inst_new_sdram_controller_0_wire_cs_n),  //        .cs_n
		.zs_dqm   (anxious_qsys_inst_new_sdram_controller_0_wire_dqm),   //        .dqm
		.zs_ras_n (anxious_qsys_inst_new_sdram_controller_0_wire_ras_n), //        .ras_n
		.zs_we_n  (anxious_qsys_inst_new_sdram_controller_0_wire_we_n)   //        .we_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) sdram_controller_0_my_partner_clk_bfm (
		.clk (sdram_controller_0_my_partner_clk_bfm_clk_clk)  // clk.clk
	);
	
	// Clock period
	localparam time CLK_PERIOD = 20ns;
	localparam time PCLK_PERIOD = 40ns;
	localparam int VSYNC_H_LINES = 1;
	localparam int VSYNC_L_LINES = 10; // Active
	localparam int HSYNC_FRONT_CYCLES = 1;
	localparam int HSYNC_ACTIVE_CYCLES = 2 * 20;
	localparam int HSYNC_BACK_CYCLES = 1;
	localparam int LINE_CYCLES = HSYNC_FRONT_CYCLES +
		HSYNC_ACTIVE_CYCLES + HSYNC_BACK_CYCLES;
	
	// Camera Signals
	logic clk_camera;
	logic [7:0] cam_din;
	logic cam_href;
	logic cam_pclk;
	logic cam_pwdn;
	logic cam_reset;
	logic cam_vsync;
	logic cam_xclk;

	logic enable_n;
	
	initial begin
		cam_pclk = 1'b0;
		camera_bfm.set_cam_pclk(cam_pclk);
	end always begin
		#(PCLK_PERIOD / 2) cam_pclk <= ~cam_pclk;
		camera_bfm.set_cam_pclk(cam_pclk);
	end

	initial begin
		clk_camera = 1'b0;
		camera_bfm.set_clk_camera(clk_camera);
	end always begin
		#(PCLK_PERIOD / 2) clk_camera <= ~clk_camera;
		camera_bfm.set_clk_camera(clk_camera);
	end

	initial begin
		cam_href = 1'b0;
		camera_bfm.set_cam_href(cam_href);
	end always begin
		#(HSYNC_FRONT_CYCLES * PCLK_PERIOD) cam_href = 1'b1;
		camera_bfm.set_cam_href(cam_href);
		#(HSYNC_ACTIVE_CYCLES * PCLK_PERIOD) cam_href = 1'b0;
		camera_bfm.set_cam_href(cam_href);
		#(HSYNC_BACK_CYCLES * PCLK_PERIOD) cam_href = 1'b0;
		camera_bfm.set_cam_href(cam_href);
	end

	initial begin
		cam_vsync = 1'b1;
		camera_bfm.set_cam_vsync(cam_vsync);
	end always begin
		#(VSYNC_H_LINES * LINE_CYCLES * PCLK_PERIOD) cam_vsync = 1'b0;
		camera_bfm.set_cam_vsync(cam_vsync);
		#(VSYNC_L_LINES * LINE_CYCLES * PCLK_PERIOD) cam_vsync = 1'b1;
		camera_bfm.set_cam_vsync(cam_vsync);
	end
	
	int row;

	initial begin
		cam_din = 2'h00;
		camera_bfm.set_cam_din(cam_din);
	end always begin
		#(VSYNC_H_LINES * LINE_CYCLES * PCLK_PERIOD) cam_din = 2'h00;
		camera_bfm.set_cam_din(cam_din);
		for (row = 0; row < 480; ++row) begin
			#(LINE_CYCLES * PCLK_PERIOD) cam_din = cam_din + 1;
			camera_bfm.set_cam_din(cam_din);
		end
	end
	
	initial begin
		camera_bfm.set_enable_n(1'b0);
		
	end

endmodule
