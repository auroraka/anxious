// mm_lock_sim_tb.v

// Generated using ACDS version 15.0 145

`timescale 1 ns / 1 ns
module mm_lock_sim_tb (
	);

	wire         mm_lock_sim_inst_clk_bfm_clk_clk;                                   // mm_lock_sim_inst_clk_bfm:clk -> [mm_lock_sim_inst:clk_clk, mm_lock_sim_inst_camera_mm_0_buffer_port_bfm:clk, mm_lock_sim_inst_camera_mm_0_conduit_bfm:clk, mm_lock_sim_inst_reset_bfm:clk, mm_lock_sim_inst_vga_composer_0_cam_buffer_bfm:clk, mm_lock_sim_inst_vga_composer_0_conduit_bfm:clk, new_sdram_controller_0_my_partner:clk]
	wire   [1:0] mm_lock_sim_inst_camera_mm_0_buffer_port_bfm_conduit_address;       // mm_lock_sim_inst_camera_mm_0_buffer_port_bfm:sig_address -> mm_lock_sim_inst:camera_mm_0_buffer_port_address
	wire   [0:0] mm_lock_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_vsync;         // mm_lock_sim_inst_camera_mm_0_conduit_bfm:sig_cam_vsync -> mm_lock_sim_inst:camera_mm_0_conduit_cam_vsync
	wire         mm_lock_sim_inst_camera_mm_0_conduit_cam_pwdn;                      // mm_lock_sim_inst:camera_mm_0_conduit_cam_pwdn -> mm_lock_sim_inst_camera_mm_0_conduit_bfm:sig_cam_pwdn
	wire   [7:0] mm_lock_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_din;           // mm_lock_sim_inst_camera_mm_0_conduit_bfm:sig_cam_din -> mm_lock_sim_inst:camera_mm_0_conduit_cam_din
	wire   [0:0] mm_lock_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_pclk;          // mm_lock_sim_inst_camera_mm_0_conduit_bfm:sig_cam_pclk -> mm_lock_sim_inst:camera_mm_0_conduit_cam_pclk
	wire   [0:0] mm_lock_sim_inst_camera_mm_0_conduit_bfm_conduit_enable_n;          // mm_lock_sim_inst_camera_mm_0_conduit_bfm:sig_enable_n -> mm_lock_sim_inst:camera_mm_0_conduit_enable_n
	wire   [0:0] mm_lock_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_href;          // mm_lock_sim_inst_camera_mm_0_conduit_bfm:sig_cam_href -> mm_lock_sim_inst:camera_mm_0_conduit_cam_href
	wire         mm_lock_sim_inst_camera_mm_0_conduit_cam_xclk;                      // mm_lock_sim_inst:camera_mm_0_conduit_cam_xclk -> mm_lock_sim_inst_camera_mm_0_conduit_bfm:sig_cam_xclk
	wire         mm_lock_sim_inst_camera_mm_0_conduit_cam_reset;                     // mm_lock_sim_inst:camera_mm_0_conduit_cam_reset -> mm_lock_sim_inst_camera_mm_0_conduit_bfm:sig_cam_reset
	wire   [0:0] mm_lock_sim_inst_camera_mm_0_conduit_bfm_conduit_clk_camera;        // mm_lock_sim_inst_camera_mm_0_conduit_bfm:sig_clk_camera -> mm_lock_sim_inst:camera_mm_0_conduit_clk_camera
	wire         mm_lock_sim_inst_new_sdram_controller_0_wire_cs_n;                  // mm_lock_sim_inst:new_sdram_controller_0_wire_cs_n -> new_sdram_controller_0_my_partner:zs_cs_n
	wire   [3:0] mm_lock_sim_inst_new_sdram_controller_0_wire_dqm;                   // mm_lock_sim_inst:new_sdram_controller_0_wire_dqm -> new_sdram_controller_0_my_partner:zs_dqm
	wire         mm_lock_sim_inst_new_sdram_controller_0_wire_cas_n;                 // mm_lock_sim_inst:new_sdram_controller_0_wire_cas_n -> new_sdram_controller_0_my_partner:zs_cas_n
	wire         mm_lock_sim_inst_new_sdram_controller_0_wire_ras_n;                 // mm_lock_sim_inst:new_sdram_controller_0_wire_ras_n -> new_sdram_controller_0_my_partner:zs_ras_n
	wire         mm_lock_sim_inst_new_sdram_controller_0_wire_we_n;                  // mm_lock_sim_inst:new_sdram_controller_0_wire_we_n -> new_sdram_controller_0_my_partner:zs_we_n
	wire  [12:0] mm_lock_sim_inst_new_sdram_controller_0_wire_addr;                  // mm_lock_sim_inst:new_sdram_controller_0_wire_addr -> new_sdram_controller_0_my_partner:zs_addr
	wire         mm_lock_sim_inst_new_sdram_controller_0_wire_cke;                   // mm_lock_sim_inst:new_sdram_controller_0_wire_cke -> new_sdram_controller_0_my_partner:zs_cke
	wire  [31:0] mm_lock_sim_inst_new_sdram_controller_0_wire_dq;                    // [] -> [mm_lock_sim_inst:new_sdram_controller_0_wire_dq, new_sdram_controller_0_my_partner:zs_dq]
	wire   [1:0] mm_lock_sim_inst_new_sdram_controller_0_wire_ba;                    // mm_lock_sim_inst:new_sdram_controller_0_wire_ba -> new_sdram_controller_0_my_partner:zs_ba
	wire   [1:0] mm_lock_sim_inst_vga_composer_0_cam_buffer_bfm_conduit_buffer_port; // mm_lock_sim_inst_vga_composer_0_cam_buffer_bfm:sig_buffer_port -> mm_lock_sim_inst:vga_composer_0_cam_buffer_buffer_port
	wire         mm_lock_sim_inst_vga_composer_0_cam_buffer_buffer_vsync;            // mm_lock_sim_inst:vga_composer_0_cam_buffer_buffer_vsync -> mm_lock_sim_inst_vga_composer_0_cam_buffer_bfm:sig_buffer_vsync
	wire         mm_lock_sim_inst_vga_composer_0_conduit_vga_clk;                    // mm_lock_sim_inst:vga_composer_0_conduit_vga_clk -> mm_lock_sim_inst_vga_composer_0_conduit_bfm:sig_vga_clk
	wire   [0:0] mm_lock_sim_inst_vga_composer_0_conduit_bfm_conduit_clk_vga;        // mm_lock_sim_inst_vga_composer_0_conduit_bfm:sig_clk_vga -> mm_lock_sim_inst:vga_composer_0_conduit_clk_vga
	wire   [7:0] mm_lock_sim_inst_vga_composer_0_conduit_vga_g;                      // mm_lock_sim_inst:vga_composer_0_conduit_vga_g -> mm_lock_sim_inst_vga_composer_0_conduit_bfm:sig_vga_g
	wire         mm_lock_sim_inst_vga_composer_0_conduit_vga_sync_n;                 // mm_lock_sim_inst:vga_composer_0_conduit_vga_sync_n -> mm_lock_sim_inst_vga_composer_0_conduit_bfm:sig_vga_sync_n
	wire         mm_lock_sim_inst_vga_composer_0_conduit_vga_vs;                     // mm_lock_sim_inst:vga_composer_0_conduit_vga_vs -> mm_lock_sim_inst_vga_composer_0_conduit_bfm:sig_vga_vs
	wire         mm_lock_sim_inst_vga_composer_0_conduit_vga_blank_n;                // mm_lock_sim_inst:vga_composer_0_conduit_vga_blank_n -> mm_lock_sim_inst_vga_composer_0_conduit_bfm:sig_vga_blank_n
	wire   [7:0] mm_lock_sim_inst_vga_composer_0_conduit_vga_b;                      // mm_lock_sim_inst:vga_composer_0_conduit_vga_b -> mm_lock_sim_inst_vga_composer_0_conduit_bfm:sig_vga_b
	wire   [7:0] mm_lock_sim_inst_vga_composer_0_conduit_vga_r;                      // mm_lock_sim_inst:vga_composer_0_conduit_vga_r -> mm_lock_sim_inst_vga_composer_0_conduit_bfm:sig_vga_r
	wire         mm_lock_sim_inst_vga_composer_0_conduit_vga_hs;                     // mm_lock_sim_inst:vga_composer_0_conduit_vga_hs -> mm_lock_sim_inst_vga_composer_0_conduit_bfm:sig_vga_hs
	wire         mm_lock_sim_inst_reset_bfm_reset_reset;                             // mm_lock_sim_inst_reset_bfm:reset -> mm_lock_sim_inst:reset_reset_n

	mm_lock_sim mm_lock_sim_inst (
		.camera_mm_0_buffer_port_address        (mm_lock_sim_inst_camera_mm_0_buffer_port_bfm_conduit_address),       //     camera_mm_0_buffer_port.address
		.camera_mm_0_conduit_clk_camera         (mm_lock_sim_inst_camera_mm_0_conduit_bfm_conduit_clk_camera),        //         camera_mm_0_conduit.clk_camera
		.camera_mm_0_conduit_enable_n           (mm_lock_sim_inst_camera_mm_0_conduit_bfm_conduit_enable_n),          //                            .enable_n
		.camera_mm_0_conduit_cam_din            (mm_lock_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_din),           //                            .cam_din
		.camera_mm_0_conduit_cam_href           (mm_lock_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_href),          //                            .cam_href
		.camera_mm_0_conduit_cam_pclk           (mm_lock_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_pclk),          //                            .cam_pclk
		.camera_mm_0_conduit_cam_pwdn           (mm_lock_sim_inst_camera_mm_0_conduit_cam_pwdn),                      //                            .cam_pwdn
		.camera_mm_0_conduit_cam_reset          (mm_lock_sim_inst_camera_mm_0_conduit_cam_reset),                     //                            .cam_reset
		.camera_mm_0_conduit_cam_vsync          (mm_lock_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_vsync),         //                            .cam_vsync
		.camera_mm_0_conduit_cam_xclk           (mm_lock_sim_inst_camera_mm_0_conduit_cam_xclk),                      //                            .cam_xclk
		.clk_clk                                (mm_lock_sim_inst_clk_bfm_clk_clk),                                   //                         clk.clk
		.new_sdram_controller_0_wire_addr       (mm_lock_sim_inst_new_sdram_controller_0_wire_addr),                  // new_sdram_controller_0_wire.addr
		.new_sdram_controller_0_wire_ba         (mm_lock_sim_inst_new_sdram_controller_0_wire_ba),                    //                            .ba
		.new_sdram_controller_0_wire_cas_n      (mm_lock_sim_inst_new_sdram_controller_0_wire_cas_n),                 //                            .cas_n
		.new_sdram_controller_0_wire_cke        (mm_lock_sim_inst_new_sdram_controller_0_wire_cke),                   //                            .cke
		.new_sdram_controller_0_wire_cs_n       (mm_lock_sim_inst_new_sdram_controller_0_wire_cs_n),                  //                            .cs_n
		.new_sdram_controller_0_wire_dq         (mm_lock_sim_inst_new_sdram_controller_0_wire_dq),                    //                            .dq
		.new_sdram_controller_0_wire_dqm        (mm_lock_sim_inst_new_sdram_controller_0_wire_dqm),                   //                            .dqm
		.new_sdram_controller_0_wire_ras_n      (mm_lock_sim_inst_new_sdram_controller_0_wire_ras_n),                 //                            .ras_n
		.new_sdram_controller_0_wire_we_n       (mm_lock_sim_inst_new_sdram_controller_0_wire_we_n),                  //                            .we_n
		.reset_reset_n                          (mm_lock_sim_inst_reset_bfm_reset_reset),                             //                       reset.reset_n
		.vga_composer_0_cam_buffer_buffer_port  (mm_lock_sim_inst_vga_composer_0_cam_buffer_bfm_conduit_buffer_port), //   vga_composer_0_cam_buffer.buffer_port
		.vga_composer_0_cam_buffer_buffer_vsync (mm_lock_sim_inst_vga_composer_0_cam_buffer_buffer_vsync),            //                            .buffer_vsync
		.vga_composer_0_conduit_vga_b           (mm_lock_sim_inst_vga_composer_0_conduit_vga_b),                      //      vga_composer_0_conduit.vga_b
		.vga_composer_0_conduit_vga_blank_n     (mm_lock_sim_inst_vga_composer_0_conduit_vga_blank_n),                //                            .vga_blank_n
		.vga_composer_0_conduit_vga_clk         (mm_lock_sim_inst_vga_composer_0_conduit_vga_clk),                    //                            .vga_clk
		.vga_composer_0_conduit_vga_g           (mm_lock_sim_inst_vga_composer_0_conduit_vga_g),                      //                            .vga_g
		.vga_composer_0_conduit_vga_hs          (mm_lock_sim_inst_vga_composer_0_conduit_vga_hs),                     //                            .vga_hs
		.vga_composer_0_conduit_vga_r           (mm_lock_sim_inst_vga_composer_0_conduit_vga_r),                      //                            .vga_r
		.vga_composer_0_conduit_vga_sync_n      (mm_lock_sim_inst_vga_composer_0_conduit_vga_sync_n),                 //                            .vga_sync_n
		.vga_composer_0_conduit_vga_vs          (mm_lock_sim_inst_vga_composer_0_conduit_vga_vs),                     //                            .vga_vs
		.vga_composer_0_conduit_clk_vga         (mm_lock_sim_inst_vga_composer_0_conduit_bfm_conduit_clk_vga)         //                            .clk_vga
	);

	altera_conduit_bfm camera_buffer_bfm (
		.clk         (mm_lock_sim_inst_clk_bfm_clk_clk),                             //     clk.clk
		.sig_address (mm_lock_sim_inst_camera_mm_0_buffer_port_bfm_conduit_address), // conduit.address
		.reset       (1'b0)                                                          // (terminated)
	);

	altera_conduit_bfm_0002 camera_bfm (
		.clk            (mm_lock_sim_inst_clk_bfm_clk_clk),                            //     clk.clk
		.sig_clk_camera (mm_lock_sim_inst_camera_mm_0_conduit_bfm_conduit_clk_camera), // conduit.clk_camera
		.sig_enable_n   (mm_lock_sim_inst_camera_mm_0_conduit_bfm_conduit_enable_n),   //        .enable_n
		.sig_cam_din    (mm_lock_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_din),    //        .cam_din
		.sig_cam_href   (mm_lock_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_href),   //        .cam_href
		.sig_cam_pclk   (mm_lock_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_pclk),   //        .cam_pclk
		.sig_cam_pwdn   (mm_lock_sim_inst_camera_mm_0_conduit_cam_pwdn),               //        .cam_pwdn
		.sig_cam_reset  (mm_lock_sim_inst_camera_mm_0_conduit_cam_reset),              //        .cam_reset
		.sig_cam_vsync  (mm_lock_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_vsync),  //        .cam_vsync
		.sig_cam_xclk   (mm_lock_sim_inst_camera_mm_0_conduit_cam_xclk),               //        .cam_xclk
		.reset          (1'b0)                                                         // (terminated)
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) mm_lock_sim_inst_clk_bfm (
		.clk (mm_lock_sim_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) mm_lock_sim_inst_reset_bfm (
		.reset (mm_lock_sim_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (mm_lock_sim_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm_0003 vga_cam_buffer_bfm (
		.clk              (mm_lock_sim_inst_clk_bfm_clk_clk),                                   //     clk.clk
		.sig_buffer_port  (mm_lock_sim_inst_vga_composer_0_cam_buffer_bfm_conduit_buffer_port), // conduit.buffer_port
		.sig_buffer_vsync (mm_lock_sim_inst_vga_composer_0_cam_buffer_buffer_vsync),            //        .buffer_vsync
		.reset            (1'b0)                                                                // (terminated)
	);

	altera_conduit_bfm_0004 vga_bfm (
		.clk             (mm_lock_sim_inst_clk_bfm_clk_clk),                            //     clk.clk
		.sig_vga_b       (mm_lock_sim_inst_vga_composer_0_conduit_vga_b),               // conduit.vga_b
		.sig_vga_blank_n (mm_lock_sim_inst_vga_composer_0_conduit_vga_blank_n),         //        .vga_blank_n
		.sig_vga_clk     (mm_lock_sim_inst_vga_composer_0_conduit_vga_clk),             //        .vga_clk
		.sig_vga_g       (mm_lock_sim_inst_vga_composer_0_conduit_vga_g),               //        .vga_g
		.sig_vga_hs      (mm_lock_sim_inst_vga_composer_0_conduit_vga_hs),              //        .vga_hs
		.sig_vga_r       (mm_lock_sim_inst_vga_composer_0_conduit_vga_r),               //        .vga_r
		.sig_vga_sync_n  (mm_lock_sim_inst_vga_composer_0_conduit_vga_sync_n),          //        .vga_sync_n
		.sig_vga_vs      (mm_lock_sim_inst_vga_composer_0_conduit_vga_vs),              //        .vga_vs
		.sig_clk_vga     (mm_lock_sim_inst_vga_composer_0_conduit_bfm_conduit_clk_vga), //        .clk_vga
		.reset           (1'b0)                                                         // (terminated)
	);

	altera_sdram_partner_module new_sdram_controller_0_my_partner (
		.clk      (mm_lock_sim_inst_clk_bfm_clk_clk),                   //     clk.clk
		.zs_dq    (mm_lock_sim_inst_new_sdram_controller_0_wire_dq),    // conduit.dq
		.zs_addr  (mm_lock_sim_inst_new_sdram_controller_0_wire_addr),  //        .addr
		.zs_ba    (mm_lock_sim_inst_new_sdram_controller_0_wire_ba),    //        .ba
		.zs_cas_n (mm_lock_sim_inst_new_sdram_controller_0_wire_cas_n), //        .cas_n
		.zs_cke   (mm_lock_sim_inst_new_sdram_controller_0_wire_cke),   //        .cke
		.zs_cs_n  (mm_lock_sim_inst_new_sdram_controller_0_wire_cs_n),  //        .cs_n
		.zs_dqm   (mm_lock_sim_inst_new_sdram_controller_0_wire_dqm),   //        .dqm
		.zs_ras_n (mm_lock_sim_inst_new_sdram_controller_0_wire_ras_n), //        .ras_n
		.zs_we_n  (mm_lock_sim_inst_new_sdram_controller_0_wire_we_n)   //        .we_n
	);
	
	// Clock period
	localparam time CLK_PERIOD = 20ns;
	localparam time PCLK_PERIOD = 40ns;
	// localparam int VSYNC_H_LINES = 3;
	// localparam int VSYNC_L_LINES = 480; // Active
	// localparam int HSYNC_FRONT_CYCLES = 144;
	// localparam int HSYNC_ACTIVE_CYCLES = 2 * 640;
	// localparam int HSYNC_BACK_CYCLES = 144;
	localparam int VSYNC_H_LINES = 1;
	localparam int VSYNC_L_LINES = 10; // Active
	localparam int HSYNC_FRONT_CYCLES = 2;
	localparam int HSYNC_ACTIVE_CYCLES = 2 * 32;
	localparam int HSYNC_BACK_CYCLES = 2;
	localparam int LINE_CYCLES = HSYNC_FRONT_CYCLES +
		HSYNC_ACTIVE_CYCLES + HSYNC_BACK_CYCLES;
	
	// Camera Signals
	logic clk_camera;
	logic [7:0] cam_din;
	logic cam_href;
	logic cam_pclk;
	logic cam_pwdn;
	logic cam_reset;
	logic cam_vsync;
	logic cam_xclk;

	logic enable_n;
	
	logic clk_vga;
	
	initial begin
		clk_vga = 1'b0;
		vga_bfm.set_clk_vga(clk_vga);
	end always begin
		#40ns clk_vga <= ~clk_vga;
		vga_bfm.set_clk_vga(clk_vga);
	end
	
	initial begin
		cam_pclk = 1'b0;
		camera_bfm.set_cam_pclk(cam_pclk);
	end always begin
		#(PCLK_PERIOD / 2) cam_pclk <= ~cam_pclk;
		camera_bfm.set_cam_pclk(cam_pclk);
	end

	initial begin
		clk_camera = 1'b0;
		camera_bfm.set_clk_camera(clk_camera);
	end always begin
		#(PCLK_PERIOD / 2) clk_camera <= ~clk_camera;
		camera_bfm.set_clk_camera(clk_camera);
	end

	initial begin
		cam_href = 1'b0;
		camera_bfm.set_cam_href(cam_href);
	end always begin
		#(HSYNC_FRONT_CYCLES * PCLK_PERIOD) cam_href = 1'b1;
		camera_bfm.set_cam_href(cam_href);
		#(HSYNC_ACTIVE_CYCLES * PCLK_PERIOD) cam_href = 1'b0;
		camera_bfm.set_cam_href(cam_href);
		#(HSYNC_BACK_CYCLES * PCLK_PERIOD) cam_href = 1'b0;
		camera_bfm.set_cam_href(cam_href);
	end

	initial begin
		cam_vsync = 1'b1;
		camera_bfm.set_cam_vsync(cam_vsync);
	end always begin
		#(VSYNC_H_LINES * LINE_CYCLES * PCLK_PERIOD) cam_vsync = 1'b0;
		camera_bfm.set_cam_vsync(cam_vsync);
		#(VSYNC_L_LINES * LINE_CYCLES * PCLK_PERIOD) cam_vsync = 1'b1;
		camera_bfm.set_cam_vsync(cam_vsync);
	end
	
	int row;

	initial begin
		cam_din = 2'h00;
		camera_bfm.set_cam_din(cam_din);
	end always begin
		#(VSYNC_H_LINES * LINE_CYCLES * PCLK_PERIOD) cam_din = 2'h00;
		camera_bfm.set_cam_din(cam_din);
		for (row = 0; row < VSYNC_L_LINES; ++row) begin
			#(LINE_CYCLES * PCLK_PERIOD) cam_din = cam_din + 1;
			camera_bfm.set_cam_din(cam_din);
		end
	end
	
	initial begin
		camera_bfm.set_enable_n(1'b0);
		camera_buffer_bfm.set_address(2'b00);
		vga_cam_buffer_bfm.set_buffer_port(2'b00);
		// wait(cam_vsync == 1'b0);
		// wait(cam_vsync == 1'b1);
		// $stop;
	end

endmodule
