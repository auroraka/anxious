// frame_buffer_sim_tb.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module frame_buffer_sim_tb (
	);

	wire        frame_buffer_sim_inst_clk_bfm_clk_clk;                            // frame_buffer_sim_inst_clk_bfm:clk -> [frame_buffer_sim_inst:clk_clk, frame_buffer_sim_inst_camera_mm_0_conduit_bfm:clk, frame_buffer_sim_inst_reset_bfm:clk, frame_buffer_sim_inst_vga_mm_0_conduit_bfm:clk]
	wire  [0:0] frame_buffer_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_vsync;  // frame_buffer_sim_inst_camera_mm_0_conduit_bfm:sig_cam_vsync -> frame_buffer_sim_inst:camera_mm_0_conduit_cam_vsync
	wire        frame_buffer_sim_inst_camera_mm_0_conduit_cam_pwdn;               // frame_buffer_sim_inst:camera_mm_0_conduit_cam_pwdn -> frame_buffer_sim_inst_camera_mm_0_conduit_bfm:sig_cam_pwdn
	wire  [7:0] frame_buffer_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_din;    // frame_buffer_sim_inst_camera_mm_0_conduit_bfm:sig_cam_din -> frame_buffer_sim_inst:camera_mm_0_conduit_cam_din
	wire  [0:0] frame_buffer_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_pclk;   // frame_buffer_sim_inst_camera_mm_0_conduit_bfm:sig_cam_pclk -> frame_buffer_sim_inst:camera_mm_0_conduit_cam_pclk
	wire  [0:0] frame_buffer_sim_inst_camera_mm_0_conduit_bfm_conduit_enable_n;   // frame_buffer_sim_inst_camera_mm_0_conduit_bfm:sig_enable_n -> frame_buffer_sim_inst:camera_mm_0_conduit_enable_n
	wire  [0:0] frame_buffer_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_href;   // frame_buffer_sim_inst_camera_mm_0_conduit_bfm:sig_cam_href -> frame_buffer_sim_inst:camera_mm_0_conduit_cam_href
	wire        frame_buffer_sim_inst_camera_mm_0_conduit_cam_xclk;               // frame_buffer_sim_inst:camera_mm_0_conduit_cam_xclk -> frame_buffer_sim_inst_camera_mm_0_conduit_bfm:sig_cam_xclk
	wire        frame_buffer_sim_inst_camera_mm_0_conduit_cam_reset;              // frame_buffer_sim_inst:camera_mm_0_conduit_cam_reset -> frame_buffer_sim_inst_camera_mm_0_conduit_bfm:sig_cam_reset
	wire  [0:0] frame_buffer_sim_inst_camera_mm_0_conduit_bfm_conduit_clk_camera; // frame_buffer_sim_inst_camera_mm_0_conduit_bfm:sig_clk_camera -> frame_buffer_sim_inst:camera_mm_0_conduit_clk_camera
	wire        frame_buffer_sim_inst_vga_mm_0_conduit_vga_clk;                   // frame_buffer_sim_inst:vga_mm_0_conduit_vga_clk -> frame_buffer_sim_inst_vga_mm_0_conduit_bfm:sig_vga_clk
	wire  [0:0] frame_buffer_sim_inst_vga_mm_0_conduit_bfm_conduit_clk_vga;       // frame_buffer_sim_inst_vga_mm_0_conduit_bfm:sig_clk_vga -> frame_buffer_sim_inst:vga_mm_0_conduit_clk_vga
	wire  [7:0] frame_buffer_sim_inst_vga_mm_0_conduit_vga_g;                     // frame_buffer_sim_inst:vga_mm_0_conduit_vga_g -> frame_buffer_sim_inst_vga_mm_0_conduit_bfm:sig_vga_g
	wire        frame_buffer_sim_inst_vga_mm_0_conduit_vga_sync_n;                // frame_buffer_sim_inst:vga_mm_0_conduit_vga_sync_n -> frame_buffer_sim_inst_vga_mm_0_conduit_bfm:sig_vga_sync_n
	wire        frame_buffer_sim_inst_vga_mm_0_conduit_vga_vs;                    // frame_buffer_sim_inst:vga_mm_0_conduit_vga_vs -> frame_buffer_sim_inst_vga_mm_0_conduit_bfm:sig_vga_vs
	wire        frame_buffer_sim_inst_vga_mm_0_conduit_vga_blank_n;               // frame_buffer_sim_inst:vga_mm_0_conduit_vga_blank_n -> frame_buffer_sim_inst_vga_mm_0_conduit_bfm:sig_vga_blank_n
	wire  [7:0] frame_buffer_sim_inst_vga_mm_0_conduit_vga_b;                     // frame_buffer_sim_inst:vga_mm_0_conduit_vga_b -> frame_buffer_sim_inst_vga_mm_0_conduit_bfm:sig_vga_b
	wire  [7:0] frame_buffer_sim_inst_vga_mm_0_conduit_vga_r;                     // frame_buffer_sim_inst:vga_mm_0_conduit_vga_r -> frame_buffer_sim_inst_vga_mm_0_conduit_bfm:sig_vga_r
	wire        frame_buffer_sim_inst_vga_mm_0_conduit_vga_hs;                    // frame_buffer_sim_inst:vga_mm_0_conduit_vga_hs -> frame_buffer_sim_inst_vga_mm_0_conduit_bfm:sig_vga_hs
	wire        frame_buffer_sim_inst_reset_bfm_reset_reset;                      // frame_buffer_sim_inst_reset_bfm:reset -> frame_buffer_sim_inst:reset_reset_n

	frame_buffer_sim frame_buffer_sim_inst (
		.camera_mm_0_conduit_clk_camera (frame_buffer_sim_inst_camera_mm_0_conduit_bfm_conduit_clk_camera), // camera_mm_0_conduit.clk_camera
		.camera_mm_0_conduit_enable_n   (frame_buffer_sim_inst_camera_mm_0_conduit_bfm_conduit_enable_n),   //                    .enable_n
		.camera_mm_0_conduit_cam_din    (frame_buffer_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_din),    //                    .cam_din
		.camera_mm_0_conduit_cam_href   (frame_buffer_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_href),   //                    .cam_href
		.camera_mm_0_conduit_cam_pclk   (frame_buffer_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_pclk),   //                    .cam_pclk
		.camera_mm_0_conduit_cam_pwdn   (frame_buffer_sim_inst_camera_mm_0_conduit_cam_pwdn),               //                    .cam_pwdn
		.camera_mm_0_conduit_cam_reset  (frame_buffer_sim_inst_camera_mm_0_conduit_cam_reset),              //                    .cam_reset
		.camera_mm_0_conduit_cam_vsync  (frame_buffer_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_vsync),  //                    .cam_vsync
		.camera_mm_0_conduit_cam_xclk   (frame_buffer_sim_inst_camera_mm_0_conduit_cam_xclk),               //                    .cam_xclk
		.clk_clk                        (frame_buffer_sim_inst_clk_bfm_clk_clk),                            //                 clk.clk
		.reset_reset_n                  (frame_buffer_sim_inst_reset_bfm_reset_reset),                      //               reset.reset_n
		.vga_mm_0_conduit_vga_b         (frame_buffer_sim_inst_vga_mm_0_conduit_vga_b),                     //    vga_mm_0_conduit.vga_b
		.vga_mm_0_conduit_vga_blank_n   (frame_buffer_sim_inst_vga_mm_0_conduit_vga_blank_n),               //                    .vga_blank_n
		.vga_mm_0_conduit_vga_clk       (frame_buffer_sim_inst_vga_mm_0_conduit_vga_clk),                   //                    .vga_clk
		.vga_mm_0_conduit_vga_g         (frame_buffer_sim_inst_vga_mm_0_conduit_vga_g),                     //                    .vga_g
		.vga_mm_0_conduit_vga_hs        (frame_buffer_sim_inst_vga_mm_0_conduit_vga_hs),                    //                    .vga_hs
		.vga_mm_0_conduit_vga_r         (frame_buffer_sim_inst_vga_mm_0_conduit_vga_r),                     //                    .vga_r
		.vga_mm_0_conduit_vga_sync_n    (frame_buffer_sim_inst_vga_mm_0_conduit_vga_sync_n),                //                    .vga_sync_n
		.vga_mm_0_conduit_vga_vs        (frame_buffer_sim_inst_vga_mm_0_conduit_vga_vs),                    //                    .vga_vs
		.vga_mm_0_conduit_clk_vga       (frame_buffer_sim_inst_vga_mm_0_conduit_bfm_conduit_clk_vga)        //                    .clk_vga
	);

	altera_conduit_bfm camera_bfm (
		.clk            (frame_buffer_sim_inst_clk_bfm_clk_clk),                            //     clk.clk
		.sig_clk_camera (frame_buffer_sim_inst_camera_mm_0_conduit_bfm_conduit_clk_camera), // conduit.clk_camera
		.sig_enable_n   (frame_buffer_sim_inst_camera_mm_0_conduit_bfm_conduit_enable_n),   //        .enable_n
		.sig_cam_din    (frame_buffer_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_din),    //        .cam_din
		.sig_cam_href   (frame_buffer_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_href),   //        .cam_href
		.sig_cam_pclk   (frame_buffer_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_pclk),   //        .cam_pclk
		.sig_cam_pwdn   (frame_buffer_sim_inst_camera_mm_0_conduit_cam_pwdn),               //        .cam_pwdn
		.sig_cam_reset  (frame_buffer_sim_inst_camera_mm_0_conduit_cam_reset),              //        .cam_reset
		.sig_cam_vsync  (frame_buffer_sim_inst_camera_mm_0_conduit_bfm_conduit_cam_vsync),  //        .cam_vsync
		.sig_cam_xclk   (frame_buffer_sim_inst_camera_mm_0_conduit_cam_xclk),               //        .cam_xclk
		.reset          (1'b0)                                                              // (terminated)
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) frame_buffer_sim_inst_clk_bfm (
		.clk (frame_buffer_sim_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) frame_buffer_sim_inst_reset_bfm (
		.reset (frame_buffer_sim_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (frame_buffer_sim_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm_0002 vga_bfm (
		.clk             (frame_buffer_sim_inst_clk_bfm_clk_clk),                      //     clk.clk
		.sig_vga_b       (frame_buffer_sim_inst_vga_mm_0_conduit_vga_b),               // conduit.vga_b
		.sig_vga_blank_n (frame_buffer_sim_inst_vga_mm_0_conduit_vga_blank_n),         //        .vga_blank_n
		.sig_vga_clk     (frame_buffer_sim_inst_vga_mm_0_conduit_vga_clk),             //        .vga_clk
		.sig_vga_g       (frame_buffer_sim_inst_vga_mm_0_conduit_vga_g),               //        .vga_g
		.sig_vga_hs      (frame_buffer_sim_inst_vga_mm_0_conduit_vga_hs),              //        .vga_hs
		.sig_vga_r       (frame_buffer_sim_inst_vga_mm_0_conduit_vga_r),               //        .vga_r
		.sig_vga_sync_n  (frame_buffer_sim_inst_vga_mm_0_conduit_vga_sync_n),          //        .vga_sync_n
		.sig_vga_vs      (frame_buffer_sim_inst_vga_mm_0_conduit_vga_vs),              //        .vga_vs
		.sig_clk_vga     (frame_buffer_sim_inst_vga_mm_0_conduit_bfm_conduit_clk_vga), //        .clk_vga
		.reset           (1'b0)                                                        // (terminated)
	);
	
	// Clock period
	localparam time CLK_PERIOD = 20ns;
	localparam time PCLK_PERIOD = 40ns;
	localparam int VSYNC_H_LINES = 3;
	localparam int VSYNC_L_LINES = 480; // Active
	localparam int HSYNC_FRONT_CYCLES = 144;
	localparam int HSYNC_ACTIVE_CYCLES = 2 * 640;
	localparam int HSYNC_BACK_CYCLES = 144;
	localparam int LINE_CYCLES = HSYNC_FRONT_CYCLES +
		HSYNC_ACTIVE_CYCLES + HSYNC_BACK_CYCLES;
	
	// Camera Signals
	logic clk_camera;
	logic [7:0] cam_din;
	logic cam_href;
	logic cam_pclk;
	logic cam_pwdn;
	logic cam_reset;
	logic cam_vsync;
	logic cam_xclk;

	logic enable_n;
	
	logic clk_vga;
	
	initial begin
		clk_vga = 1'b0;
		vga_bfm.set_clk_vga(clk_vga);
	end always begin
		#40ns clk_vga <= ~clk_vga;
		vga_bfm.set_clk_vga(clk_vga);
	end
	
	initial begin
		cam_pclk = 1'b0;
		camera_bfm.set_cam_pclk(cam_pclk);
	end always begin
		#(PCLK_PERIOD / 2) cam_pclk <= ~cam_pclk;
		camera_bfm.set_cam_pclk(cam_pclk);
	end

	initial begin
		clk_camera = 1'b0;
		camera_bfm.set_clk_camera(clk_camera);
	end always begin
		#(PCLK_PERIOD / 2) clk_camera <= ~clk_camera;
		camera_bfm.set_clk_camera(clk_camera);
	end

	initial begin
		cam_href = 1'b0;
		camera_bfm.set_cam_href(cam_href);
	end always begin
		#(HSYNC_FRONT_CYCLES * PCLK_PERIOD) cam_href = 1'b1;
		camera_bfm.set_cam_href(cam_href);
		#(HSYNC_ACTIVE_CYCLES * PCLK_PERIOD) cam_href = 1'b0;
		camera_bfm.set_cam_href(cam_href);
		#(HSYNC_BACK_CYCLES * PCLK_PERIOD) cam_href = 1'b0;
		camera_bfm.set_cam_href(cam_href);
	end

	initial begin
		cam_vsync = 1'b1;
		camera_bfm.set_cam_vsync(cam_vsync);
	end always begin
		#(VSYNC_H_LINES * LINE_CYCLES * PCLK_PERIOD) cam_vsync = 1'b0;
		camera_bfm.set_cam_vsync(cam_vsync);
		#(VSYNC_L_LINES * LINE_CYCLES * PCLK_PERIOD) cam_vsync = 1'b1;
		camera_bfm.set_cam_vsync(cam_vsync);
	end
	
	int row;

	initial begin
		cam_din = 2'h00;
		camera_bfm.set_cam_din(cam_din);
	end always begin
		#(VSYNC_H_LINES * LINE_CYCLES * PCLK_PERIOD) cam_din = 2'h00;
		camera_bfm.set_cam_din(cam_din);
		for (row = 0; row < VSYNC_L_LINES; ++row) begin
			#(LINE_CYCLES * PCLK_PERIOD) cam_din = cam_din + 1;
			camera_bfm.set_cam_din(cam_din);
		end
	end
	
	initial begin
		camera_bfm.set_enable_n(1'b0);
		wait(cam_vsync == 1'b0);
		wait(cam_vsync == 1'b1);
		$stop;
	end

endmodule
